package types;

    

endpackage