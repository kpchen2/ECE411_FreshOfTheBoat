// module top_tb;

//     timeunit 1ps;
//     timeprecision 1ps;

//     int clock_half_period_ps;
//     initial begin
//         $value$plusargs("CLOCK_PERIOD_PS_ECE411=%d", clock_half_period_ps);
//         clock_half_period_ps = clock_half_period_ps / 2;
//     end

//     bit clk;
//     always #(clock_half_period_ps) clk = ~clk;

//     bit rst;

//     int timeout = 10000000; // in cycles, change according to your needs

//     mem_itf_banked mem_itf(.*);
//     dram_w_burst_frfcfs_controller mem(.itf(mem_itf));

//     mon_itf #(.CHANNELS(8)) mon_itf(.*);
//     monitor #(.CHANNELS(8)) monitor(.itf(mon_itf));

//     cpu dut(
//         .clk            (clk),
//         .rst            (rst),

//         .bmem_addr  (mem_itf.addr  ),
//         .bmem_read  (mem_itf.read  ),
//         .bmem_write (mem_itf.write ),
//         .bmem_wdata (mem_itf.wdata ),
//         .bmem_ready (mem_itf.ready ),
//         .bmem_raddr (mem_itf.raddr ),
//         .bmem_rdata (mem_itf.rdata ),
//         .bmem_rvalid(mem_itf.rvalid)
//     );

//     `include "rvfi_reference.svh"

//     initial begin
//         $fsdbDumpfile("dump.fsdb");
//         $fsdbDumpvars(0, "+all");
//         rst = 1'b1;
//         repeat (2) @(posedge clk);
//         rst <= 1'b0;
//     end

//     always @(posedge clk) begin
//         for (int unsigned i=0; i < 8; ++i) begin
//             if (mon_itf.halt[i]) begin
//                 $finish;
//             end
//         end
//         if (timeout == 0) begin
//             $error("TB Error: Timed out");
//             $finish;
//         end
//         if (mon_itf.error != 0) begin
//             repeat (5) @(posedge clk);
//             $finish;
//         end
//         if (mem_itf.error != 0) begin
//             repeat (5) @(posedge clk);
//             $finish;
//         end
//         timeout <= timeout - 1;
//     end

// endmodule
